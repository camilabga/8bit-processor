library verilog;
use verilog.vl_types.all;
entity phasePWM_mode_vlg_vec_tst is
end phasePWM_mode_vlg_vec_tst;
