library verilog;
use verilog.vl_types.all;
entity shr_8bits_vlg_vec_tst is
end shr_8bits_vlg_vec_tst;
