library verilog;
use verilog.vl_types.all;
entity mult_8bits_vlg_vec_tst is
end mult_8bits_vlg_vec_tst;
