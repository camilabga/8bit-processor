library verilog;
use verilog.vl_types.all;
entity banco_ABCD_vlg_vec_tst is
end banco_ABCD_vlg_vec_tst;
