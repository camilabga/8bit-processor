library verilog;
use verilog.vl_types.all;
entity seletor_moeda_vlg_vec_tst is
end seletor_moeda_vlg_vec_tst;
