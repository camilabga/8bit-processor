library verilog;
use verilog.vl_types.all;
entity lab06_vlg_vec_tst is
end lab06_vlg_vec_tst;
