library verilog;
use verilog.vl_types.all;
entity lab03_vlg_vec_tst is
end lab03_vlg_vec_tst;
