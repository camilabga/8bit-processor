library verilog;
use verilog.vl_types.all;
entity lab04_vlg_vec_tst is
end lab04_vlg_vec_tst;
