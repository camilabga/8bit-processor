library verilog;
use verilog.vl_types.all;
entity SD07_vlg_vec_tst is
end SD07_vlg_vec_tst;
