library verilog;
use verilog.vl_types.all;
entity fastPWM_mode_vlg_vec_tst is
end fastPWM_mode_vlg_vec_tst;
