library verilog;
use verilog.vl_types.all;
entity select_mux_rom_vlg_vec_tst is
end select_mux_rom_vlg_vec_tst;
