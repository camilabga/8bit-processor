library verilog;
use verilog.vl_types.all;
entity ctc_mode_vlg_vec_tst is
end ctc_mode_vlg_vec_tst;
