library verilog;
use verilog.vl_types.all;
entity contador16bits_vlg_vec_tst is
end contador16bits_vlg_vec_tst;
