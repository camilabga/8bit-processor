library verilog;
use verilog.vl_types.all;
entity subtrator8bits_vlg_vec_tst is
end subtrator8bits_vlg_vec_tst;
