library verilog;
use verilog.vl_types.all;
entity processador_perifericos_timer_spi_vlg_vec_tst is
end processador_perifericos_timer_spi_vlg_vec_tst;
