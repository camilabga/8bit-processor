library verilog;
use verilog.vl_types.all;
entity shl_8bits_vlg_vec_tst is
end shl_8bits_vlg_vec_tst;
