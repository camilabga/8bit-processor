library verilog;
use verilog.vl_types.all;
entity maquina_troco_vlg_vec_tst is
end maquina_troco_vlg_vec_tst;
