library verilog;
use verilog.vl_types.all;
entity timer_vlg_check_tst is
    port(
        timer0          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end timer_vlg_check_tst;
