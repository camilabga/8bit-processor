library verilog;
use verilog.vl_types.all;
entity lab01_vlg_vec_tst is
end lab01_vlg_vec_tst;
