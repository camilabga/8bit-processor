library verilog;
use verilog.vl_types.all;
entity SPI_SD_vlg_vec_tst is
end SPI_SD_vlg_vec_tst;
