library verilog;
use verilog.vl_types.all;
entity normal_mode_vlg_vec_tst is
end normal_mode_vlg_vec_tst;
