library verilog;
use verilog.vl_types.all;
entity normal_mode_vlg_check_tst is
    port(
        timer           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end normal_mode_vlg_check_tst;
