library verilog;
use verilog.vl_types.all;
entity lab05_vlg_vec_tst is
end lab05_vlg_vec_tst;
