library verilog;
use verilog.vl_types.all;
entity lab02_vlg_vec_tst is
end lab02_vlg_vec_tst;
